library verilog;
use verilog.vl_types.all;
entity sistemaComputacional_vlg_vec_tst is
end sistemaComputacional_vlg_vec_tst;
