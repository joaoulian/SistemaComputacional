module memoriaDeInstrucoes (endereco,
									 instrucao,
									 clock);
	
	//Entradas
	input [31:0] 	endereco;
	input clock;
	
	//Saidas
	output [31:0] 	instrucao;
	
	//Variaveis locais
	reg [31:0] memoriaDeInstrucoes [130:0];
	
	integer PrimeiroClock = 0;
		
	always @ (posedge clock) begin
		if (PrimeiroClock == 0) begin
			memoriaDeInstrucoes[1] = {5'd16, 27'd39};
			memoriaDeInstrucoes[2] = {5'd25, 5'd1, 22'd0};
			memoriaDeInstrucoes[3] = {5'd24, 5'd1, 22'd6};
			memoriaDeInstrucoes[4] = {5'd25, 5'd1, 22'd1};
			memoriaDeInstrucoes[5] = {5'd24, 5'd1, 22'd7};
			memoriaDeInstrucoes[6] = {5'd25, 5'd1, 22'd0};
			memoriaDeInstrucoes[7] = {5'd24, 5'd1, 22'd4};
			memoriaDeInstrucoes[8] = {5'd23, 5'd1, 22'd4};
			memoriaDeInstrucoes[9] = {5'd23, 5'd2, 22'd3};
			memoriaDeInstrucoes[10] = {5'd30, 5'd1, 5'd2, 5'd3, 12'dx};
			memoriaDeInstrucoes[11] = {5'd25, 5'd0, 22'd0};
			memoriaDeInstrucoes[12] = {5'd12, 5'd3, 5'd0, 17'd36};
			memoriaDeInstrucoes[13] = {5'd23, 5'd1, 22'd4};
			memoriaDeInstrucoes[14] = {5'd25, 5'd2, 22'd1};
			memoriaDeInstrucoes[15] = {5'd30, 5'd1, 5'd2, 5'd3, 12'dx};
			memoriaDeInstrucoes[16] = {5'd25, 5'd0, 22'd0};
			memoriaDeInstrucoes[17] = {5'd12, 5'd3, 5'd0, 17'd21};
			memoriaDeInstrucoes[18] = {5'd23, 5'd1, 22'd4};
			memoriaDeInstrucoes[19] = {5'd24, 5'd1, 22'd5};
			memoriaDeInstrucoes[20] = {5'd16, 27'd30};
			memoriaDeInstrucoes[21] = {5'd23, 5'd1, 22'd6};
			memoriaDeInstrucoes[22] = {5'd23, 5'd2, 22'd7};
			memoriaDeInstrucoes[23] = {5'd1, 5'd1, 5'd2, 5'd3, 12'dx};
			memoriaDeInstrucoes[24] = {5'd22, 5'd3, 5'd4, 17'd0};
			memoriaDeInstrucoes[25] = {5'd24, 5'd4, 22'd5};
			memoriaDeInstrucoes[26] = {5'd23, 5'd1, 22'd7};
			memoriaDeInstrucoes[27] = {5'd24, 5'd1, 22'd6};
			memoriaDeInstrucoes[28] = {5'd23, 5'd1, 22'd5};
			memoriaDeInstrucoes[29] = {5'd24, 5'd1, 22'd7};
			memoriaDeInstrucoes[30] = {5'd23, 5'd1, 22'd4};
			memoriaDeInstrucoes[31] = {5'd25, 5'd2, 22'd1};
			memoriaDeInstrucoes[32] = {5'd1, 5'd1, 5'd2, 5'd3, 12'dx};
			memoriaDeInstrucoes[33] = {5'd22, 5'd3, 5'd4, 17'd0};
			memoriaDeInstrucoes[34] = {5'd24, 5'd4, 22'd4};
			memoriaDeInstrucoes[35] = {5'd16, 27'd8};
			memoriaDeInstrucoes[36] = {5'd23, 5'd30, 22'd5};
			memoriaDeInstrucoes[37] = {5'd23, 5'd32, 22'd2};
			memoriaDeInstrucoes[38] = {5'd27, 5'd32, 22'd0};
			memoriaDeInstrucoes[39] = {5'd19, 5'd4, 22'd0};
			memoriaDeInstrucoes[40] = {5'd24, 5'd4, 22'd9};
			memoriaDeInstrucoes[41] = {5'd23, 5'd1, 22'd9};
			memoriaDeInstrucoes[42] = {5'd24, 5'd1, 22'd3};
			memoriaDeInstrucoes[43] = {5'd25, 5'd32, 22'd46};
			memoriaDeInstrucoes[44] = {5'd24, 5'd32, 22'd2};
			memoriaDeInstrucoes[45] = {5'd16, 27'd2};
			memoriaDeInstrucoes[46] = {5'd24, 5'd30, 22'd10};
			memoriaDeInstrucoes[47] = {5'd23, 5'd1, 22'd10};
			memoriaDeInstrucoes[48] = {5'd20, 5'd1, 22'd0};
			memoriaDeInstrucoes[49] = {5'd18, 27'dx};
			PrimeiroClock <= 1;
		end
	end
		
	assign instrucao = memoriaDeInstrucoes[endereco[9:0]];
	
endmodule 